----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:12:15 09/20/2024 
-- Design Name: 
-- Module Name:    my_MULTIPLIER1BIT - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity my_MULTIPLIER1BIT is
    Port ( A : in  STD_LOGIC_VECTOR;
           B : in  STD_LOGIC;
           Y : out  STD_LOGIC);
end my_MULTIPLIER1BIT;

architecture Behavioral of my_MULTIPLIER1BIT is

begin


end Behavioral;

