`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:19:07 09/20/2024 
// Design Name: 
// Module Name:    my_MULTIPLIER4BITS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module my_MULTIPLIER4BITS(
    input [3:0] A,
    input [3:0] B,
    output [3:0] Y
    );


endmodule
